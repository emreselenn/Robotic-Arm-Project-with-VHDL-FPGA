library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--------------------------------------------------------------------------------
-- 10x10 bitmap ROM VHDL_Module of English characters and digits.
-- Made by Yunus Emre SELEN
-- 22.12.2024
--------------------------------------------------------------------------------
entity RAM is
    Port (
        address : in  std_logic_vector(8 downto 0); -- 9-bit adresleme (512 satr)
        data    : out std_logic_vector(9 downto 0)
    );
end RAM;
architecture Behavioral of RAM is
    type rom_type is array (0 to 511) of std_logic_vector(9 downto 0);
    constant ROM_DATA : rom_type := (
        
		0  	=> "0000000000", -- 'A' 
        1 	=> "0011111100",  
        2 	=> "0100000010",  
        3  	=> "0100000010",  
        4 	=> "0111111110",  
        5  	=> "0100000010",  
        6 	=> "0100000010",  
        7 	=> "0100000010",  
        8  	=> "0100000010",
		9	=> "0000000000",
		
		10	=> "0000000000", -- 'B' 
        11 	=> "0011111110", 
        12 	=> "0100000010", 
        13 	=> "0100000010", 
        14 	=> "0011111110", 
        15 	=> "0100000010", 
        16 	=> "0100000010", 
        17 	=> "0100000010", 
        18 	=> "0011111110",
		19	=> "0000000000",
		
		20	=> "0000000000", -- 'C'   
		21  => "0011111100",  
        22  => "0100000010",  
        23  => "0000000010",  
        24  => "0000000010",  
        25  => "0000000010",  
        26  => "0000000010",  
        27  => "0100000010",  
        28  => "0011111100",
		29	=> "0000000000",
		
		30 	=> "0000000000", -- 'D' 
        31 	=> "0001111110", 
        32	=> "0010000010", 
        33 	=> "0100000010", 
        34	=> "0100000010", 
        35 	=> "0100000010", 
        36 	=> "0100000010", 
        37 	=> "0010000010", 
        38 	=> "0001111110", 
		39	=> "0000000000",
		
		40	=> "0000000000", -- 'E' 
        41 	=> "0111111110",
        42 	=> "0000000010",
        43 	=> "0000000010",
        44 	=> "0011111110",
        45 	=> "0000000010",
        46 	=> "0000000010",
        47 	=> "0000000010",
        48 	=> "0111111110",
		49	=> "0000000000",
		
		50  => "0000000000", -- 'F' 
        51 	=> "0111111110",
        52 	=> "0000000010",
        53 	=> "0000000010",
        54 	=> "0011111110",
        55 	=> "0000000010",
        56 	=> "0000000010",
        57 	=> "0000000010",
        58 	=> "0000000010",
		59	=> "0000000000",
		
		60	=> "0000000000", -- 'G'
		  61  => "0011111110",
        62 	=> "0100000010",
        63 	=> "0000000010",
        64 	=> "0011110010",
        65 	=> "0010000010",
        66 	=> "0100000010",
        67 	=> "0100000010",
        68 	=> "0011111100",
		69	=> "0000000000",
		
		70	=> "0000000000", -- 'H' 
        71 	=> "0100000010",
        72 	=> "0100000010",
        73 	=> "0100000010",
        74 	=> "0111111110",
        75 	=> "0100000010",
        76 	=> "0100000010",
        77 	=> "0100000010",
        78 	=> "0100000010",
		79	=> "0000000000",
		
		80	=> "0000000000", -- 'I' 
        81 	=> "0111111110",
        82 	=> "0000110000",
        83 	=> "0000110000",
        84 	=> "0000110000",
        85 	=> "0000110000",
        86 	=> "0000110000",
        87 	=> "0000110000",
        88 	=> "0111111110",
		89	=> "0000000000",	
		
		90	=> "0000000000", -- 'J' 
        91 	=> "0011110000",
        92 	=> "0100000000",
        93 	=> "0100000000",
        94 	=> "0100000000",
        95 	=> "0100000010",
        96 	=> "0100000010",
        97 	=> "0100000010",
        98 	=> "0011111100",
		99	=> "0000000000", 
		
		100	=> "0000000000", -- 'K' 
        101	=> "0100000110",
        102 => "0001000110",
        103 => "0000100110",
        104 => "0000010110",
        105 => "0000100110",
        106 => "0001000110",
        107 => "0010000110",
        108 => "0100000110",
		109	=> "0000000000",  
		
		110	=> "0000000000", -- 'L' 
        111	=> "0000000010",
        112	=> "0000000010",
        113	=> "0000000010",
        114	=> "0000000010",
        115	=> "0000000010",
        116	=> "0000000010",
        117	=> "0000000010",
        118	=> "0111111110",
		119	=> "0000000000",
		
		120	=> "0000000000", -- 'M' 
        121	=> "0100000010",
        122	=> "0011000110",
        123	=> "0010101010",
        124	=> "0010010010",
        125	=> "0010000010",
        126	=> "0010000010",
        127	=> "0010000010",
        128	=> "0010000010",
		129	=> "0000000000",  
		
		130	=> "0000000000", -- 'N' 
        131	=> "0100000010",
        132	=> "0100000110",
        133	=> "0100001010",
        134	=> "0100010010",
        135	=> "0100100010",
        136	=> "0101000010",
        137	=> "0110000010",
        138	=> "0100000010",
		139	=> "0000000000", 
		
		140	=> "0000000000", -- 'O' 
        141	=> "0011111100",
        142	=> "0100000010",
        143	=> "0100000010",
        144	=> "0100000010",
        145	=> "0100000010",
        146	=> "0100000010",
        147	=> "0100000010",
        148	=> "0011111100",
		149	=> "0000000000",
		
		150	=> "0000000000", -- 'P' 
        151	=> "0011111100",
        152	=> "0100000010",
        153	=> "0100000010",
        154	=> "0100000010",
        155	=> "0011111100",
        156	=> "0000000010",
        157	=> "0000000010",
        158	=> "0000000010",
		159	=> "0000000000", 
		
		160	=> "0000000000", --	'Q' 
        161	=> "0011111100",
        162	=> "0100000010",
        163	=> "0100000010",
        164	=> "0100000010",
        165	=> "0100000010",
        166	=> "0100100010",
        167	=> "0101000010",
        168	=> "0110111100",
		169	=> "0000000000", 
		
		170	=> "0000000000", --	'R' 
        171	=> "0011111100",
        172	=> "0100000010",
        173	=> "0100000010",
        174	=> "0100000010",
        175	=> "0011111100",
        176	=> "0001000010",
        177	=> "0010000010",
        178	=> "0100000010",
		179	=> "0000000000",  
		
		180	=> "0000000000", -- 'S' 
        181	=> "0111111100",
        182	=> "0000000010",
        183	=> "0000000010",
        184	=> "0011111100",
        185	=> "0100000000",
        186	=> "0100000000",
        187	=> "0100000000",
        188	=> "0011111110",
		189	=> "0000000000",
		
		190	=> "0000000000", --	'T' 
        191	=> "0111111110",
        192	=> "0000110000",
        193	=> "0000110000",
        194	=> "0000110000",
        195	=> "0000110000",
        196	=> "0000110000",
        197 => "0000110000",
        198	=> "0000110000",
		199	=> "0000000000",	
		
		200	=> "0000000000", -- 'U' 
		201	=> "0100000010",
		202	=> "0100000010",
		203	=> "0100000010",
		204	=> "0100000010",
		205	=> "0100000010",
		206	=> "0100000010",
		207	=> "0100000010",
		208	=> "0011111100",
		209	=> "0000000000",   
		
		210	=> "0000000000",  -- 'V' 
		211	=> "0100000010",
		212	=> "0100000010",
		213	=> "0100000010",
		214	=> "0100000010",
		215	=> "0010000100",
		216	=> "0010000100",
		217	=> "0001111000",
		218	=> "0000110000",
		219	=> "0000000000",   
		
		220	=> "0000000000", -- 'W' 
		221	=> "0100000010",
		222	=> "0100000010",
		223	=> "0100000010",
		224	=> "0100100010",
		225	=> "0101010010",
		226	=> "0101010010",
		227	=> "0110001110",
		228	=> "0100001100",
		229	=> "0000000000", 
		
		230	=> "0000000000", -- 'X' 
		231	=> "0100000010",
		232	=> "0010000100",
		233	=> "0001001000",
		234	=> "0000110000",
		235	=> "0000110000",
		236	=> "0001001000",
		237	=> "0010000100",
		238	=> "0100000010",
		239	=> "0000000000",  
		
		240	=> "0000000000", -- 'Y' 
		241	=> "0100000010",
		242	=> "0010000100",
		243	=> "0001001000",
		244	=> "0000110000",
		245	=> "0000100000",
		246	=> "0000100000",
		247	=> "0000100000",
		248	=> "0000100000",
		249	=> "0000000000",   
		
		250	=> "0000000000", -- 'Z' 
		251	=> "0111111110",
		252	=> "0100000000",
		253	=> "0010000000",
		254	=> "0001000000",
		255	=> "0000100000",
		256	=> "0000010000",
		257	=> "0000001000",
		258	=> "0111111110",
		259	=> "0000000000",	
		
		260	=> "0000000000",  -- '0' 
		261	=> "0011111100",
		262	=> "0100000010",
		263	=> "0100000010",
		264	=> "0100000010",
		265	=> "0100000010",
		266	=> "0100000010",
		267	=> "0100000010",
		268	=> "0011111100",
		269	=> "0000000000",   
		
		270	=> "0000000000", -- '1' 
		271	=> "0000100000",
		272	=> "0000110000",
		273	=> "0000101000",
		274	=> "0000100000",
		275	=> "0000100000",
		276	=> "0000100000",
		277	=> "0000100000",
		278	=> "0011111100",
		279	=> "0000000000",	
		
		280	=> "0000000000",  -- '2' 
		281	=> "0011111100",
		282	=> "0100000010",
		283	=> "0100000000",
		284	=> "0011000000",
		285	=> "0000110000",
		286	=> "0000011000",
		287	=> "0000001100",
		288	=> "0111111110",
		289	=> "0000000000", 
		
		290	=> "0000000000", -- '3' 
		291	=> "0111111110",
		292	=> "0100000000",
		293	=> "0100000000",
		294	=> "0111111100",
		295	=> "0100000000",
		296	=> "0100000000",
		297	=> "0100000000",
		298	=> "0111111110",
		299	=> "0000000000",  
		
		300	=> "0000000000", -- '4' 
		301	=> "0010000010",
		302	=> "0010000010",
		303	=> "0010000010",
		304	=> "0010000010",
		305	=> "0111111110",
		306	=> "0010000000",
		307	=> "0010000000",
		308	=> "0010000000",
		309	=> "0000000000", 
		
		310	=> "0000000000", -- '5' 
		311	=> "0111111110",
		312	=> "0000000010",
		313	=> "0000000010",
		314	=> "0111111110",
		315	=> "0100000000",
		316	=> "0100000000",
		317	=> "0100000000",
		318	=> "0011111100",
		319	=> "0000000000", 
		
		320	=> "0000000000", -- '6' 
		321	=> "0011111100",
		322	=> "0100000010",
		323	=> "0000000010",
		324	=> "0000000010",
		325	=> "0011111100",
		326	=> "0100000010",
		327	=> "0100000010",
		328	=> "0011111100",
		329	=> "0000000000",  
		
		330	=> "0000000000", -- '7' 
		331	=> "0111111110",
		332	=> "0100000000",
		333	=> "0010000000",
		334	=> "0001000000",
		335	=> "0000100000",
		336	=> "0000010000",
		337	=> "0000001000",
		338	=> "0000001000",
		339	=> "0000000000",   
		
		340	=> "0000000000", -- '8' 
		341	=> "0011111100",
		342	=> "0100000010",
		343	=> "0100000010",
		344	=> "0011111100",
		345	=> "0100000010",
		346	=> "0100000010",
		347	=> "0100000010",
		348	=> "0011111100",
		349	=> "0000000000",   
		
		350	=> "0000000000",  -- '9' 
		351	=> "0011111100",
		352	=> "0100000010",
		353	=> "0100000010",
		354	=> "0111111110",
		355	=> "0100000000",
		356	=> "0100000000",
		357	=> "0100000010",
		358	=> "0011111100",
		359	=> "0000000000",
		
		360	=> "0000000000",  -- '|' 
		361	=> "0000110000",  -- 'v'
		362	=> "0000110000",
		363	=> "0000110000",
		364	=> "0100110010",
		365	=> "0100110010",
		366	=> "0010110100",
		367	=> "0001111000",
		368	=> "0000110000",
		369	=> "0000000000",
		
		370	=> "0000000000",  -- 'x'
		371	=> "0000000000",  
		372	=> "0000000000",
		373	=> "0010000100",
		374	=> "0001001000",
		375	=> "0000110000",
		376	=> "0000110000",
		377	=> "0001001000",
		378	=> "0010000100",
		379	=> "0000000000",
		
		380	=> "0000000000",  -- 'heart'
		381	=> "0000000000",  
		382	=> "0011001100",
		383	=> "0111111110",
		384	=> "0111111110",
		385	=> "0111111110",
		386	=> "0011111100",
		387	=> "0001111000",
		388	=> "0000110000",
		389	=> "0000000000",
		
		390	=> "0000000000",  -- '/'
		391	=> "0000000010",  
		392	=> "0000000100",
		393	=> "0000001000",
		394	=> "0000010000",
		395	=> "0000100000",
		396	=> "0001000000",
		397	=> "0010000000",
		398	=> "0100000000",
		399	=> "0000000000",
         
		others => "0000000000"
		  
    );
begin
    process(address)
    begin
        data <= ROM_DATA(to_integer(unsigned(address)));
    end process;
end Behavioral;